module boid_accelerator(
	input
);

endmodule