module d_reg
	#(
		parameter d_width = 32,
		parameter d_res_v = 0
	)(
	input logic 	clk,
	input logic 	reset,
	input logic 	[d_width-1:0] d,
	output logic 	[d_width-1:0] q
	);
	
	always @(posedge clk) begin
		if (reset) begin
			q <= d_res_v;
		end else begin
			q <= d;
		end
	end
	
endmodule

module fix15_mul(
	input logic signed 	[31:0] a, b,
	output logic signed	[31:0] q
	);
	
	logic signed [63:0] temp;
	assign temp = a * b;
	assign q = temp >>> 15;
	
endmodule

module amax_bmin(
	input logic 	[31:0] a, b,
	output logic	[31:0] q
	);
	
	logic signed [31:0] 	a_temp, 	b_temp,
								a_out,	b_out;
	
	logic signed [31:0] alpha, beta;
	
	fix15_mul a_mul(
		.a(a),
		.b(32'hffff0000),
		.q(a_out)
		);
		
	fix15_mul b_mul(
		.a(32'hffff0000),
		.b(b),
		.q(b_out)
		);
	
	
	
	//absolute value
	always_comb begin
		if (a[31] == 1) begin
			a_temp = a_out + (32'b1);
		end else begin
			a_temp = a;
		end
		
		if (b[31] == 1) begin
			b_temp = b_out + (32'b1);
		end else begin
			b_temp = b;
		end		
		
		if (a > b) begin
			alpha = a_temp;
			beta = b_temp;
		end else begin
			alpha = b_temp;
			beta = a_temp;
		end
		
		q = alpha + (beta >>> 1);
		
	end
	
	
endmodule

// fall_edge_detector will pulse 1 cycle high when a falling edge is recorded (with 1 cycle delay)

module fall_edge_detector(
  input  logic clk, signal,
  output logic q
);

  logic signalPrev;

  always_ff @(posedge clk) begin
    signalPrev <= signal;
    q       <= (!signal && signalPrev);
  end

endmodule

// zero_pad_fix15 will sign extend the variable on fix_in to 32 bits, with 
// compile-time defined parameters to determine how it should be interpreted.
// on a [total_bit_width - 1:0] register, the variable to be sign extended
// will be on bits [ (16 + fix_whole_bit_width + lsb_offset) : lsb_offset]
// and the sign will be on bit 16 + fix_whole_bit_width + lsb_offset.
// Requirement: total_bit_width, as defined, must be equal to or greater than 
// 16 + fix_whole_bit_width + lsb_offset.

module zero_pad_fix15
#(	
	parameter fix_whole_bit_width = 16,
	parameter total_bit_width		= 32
)
(	
	input 	[fix_whole_bit_width - 1:0] fix_in,
	output	[31:0]						fix_out
);
	localparam input_fix_bit_width = fix_whole_bit_width;
	assign fix_out = 
		{{(33 - input_fix_bit_width){fix_in[input_fix_bit_width - 1]}}, fix_in[input_fix_bit_width - 2:0] };

endmodule

module lut_32_divider
(	
	input logic [5:0] lut_sel,
	output logic signed[31:0] div_val
);
	// Lookup table for values of lut_sel mapping to 1/lut_sel for values
	// from 1 to 31, and returning 0 for lut_sel = 0. This will lead to
	// the centering and matching factors being zeroed out if no neighboring boids are detected.
	
	always @(*) begin
		case(lut_sel)
			0: 	div_val = 32'b0;
			1: 	div_val = 32'd1 << 16;
			2: 	div_val = 32'h00004000;
			3: 	div_val = 32'h00002aaa;
			4: 	div_val = 32'h00002000;
			5: 	div_val = 32'h00001999;
			6: 	div_val = 32'h00001555;
			7: 	div_val = 32'h00001249;
			8: 	div_val = 32'h00001000;
			9: 	div_val = 32'h00000e38;
			10: 	div_val = 32'h00000ccc;
			11: 	div_val = 32'h00000ba2;
			12: 	div_val = 32'h00000aaa;
			13: 	div_val = 32'h000009d8;
			14: 	div_val = 32'h00000924;
			15: 	div_val = 32'h00000888;
			16: 	div_val = 32'h00000800;
			17: 	div_val = 32'h00000787;
			18: 	div_val = 32'h0000071c;
			19: 	div_val = 32'h000006bc;
			20: 	div_val = 32'h00000666;
			21: 	div_val = 32'h00000618;
			22: 	div_val = 32'h000005d1;
			23: 	div_val = 32'h00000590;
			24: 	div_val = 32'h00000555;
			25: 	div_val = 32'h0000051e;
			26: 	div_val = 32'h000004ec;
			27: 	div_val = 32'h000004bd;
			28: 	div_val = 32'h00000492;
			29: 	div_val = 32'h00000469;
			30: 	div_val = 32'h00000444;
			31: 	div_val = 32'h00000421;
			default: div_val = 32'b0;
		endcase
	end

endmodule

module lut_128_divider
(	
	input logic [7:0] lut_sel,
	output logic signed[31:0] div_val
);
	always @(*) begin
		case(lut_sel)
			0: 	div_val = 32'b0;
			1: 	div_val = 32'd1 << 16;
			2: 	div_val = 32'h00004000;
			3: 	div_val = 32'h00002aaa;
			4: 	div_val = 32'h00002000;
			5: 	div_val = 32'h00001999;
			6: 	div_val = 32'h00001555;
			7: 	div_val = 32'h00001249;
			8: 	div_val = 32'h00001000;
			9: 	div_val = 32'h00000e38;
			10: 	div_val = 32'h00000ccc;
			11: 	div_val = 32'h00000ba2;
			12: 	div_val = 32'h00000aaa;
			13: 	div_val = 32'h000009d8;
			14: 	div_val = 32'h00000924;
			15: 	div_val = 32'h00000888;
			16: 	div_val = 32'h00000800;
			17: 	div_val = 32'h00000787;
			18: 	div_val = 32'h0000071c;
			19: 	div_val = 32'h000006bc;
			20: 	div_val = 32'h00000666;
			21: 	div_val = 32'h00000618;
			22: 	div_val = 32'h000005d1;
			23: 	div_val = 32'h00000590;
			24: 	div_val = 32'h00000555;
			25: 	div_val = 32'h0000051e;
			26: 	div_val = 32'h000004ec;
			27: 	div_val = 32'h000004bd;
			28: 	div_val = 32'h00000492;
			29: 	div_val = 32'h00000469;
			30: 	div_val = 32'h00000444;
			31: 	div_val = 32'h00000421;
			32: 	div_val = 32'h00000400;
			33: 	div_val = 32'h000003e0;
			34: 	div_val = 32'h000003c3;
			35: 	div_val = 32'h000003a8;
			36: 	div_val = 32'h0000038e;
			37: 	div_val = 32'h00000375;
			38: 	div_val = 32'h0000035e;
			39: 	div_val = 32'h00000348;
			40: 	div_val = 32'h00000333;
			41: 	div_val = 32'h0000031f;
			42: 	div_val = 32'h0000030c;
			43: 	div_val = 32'h000002fa;
			44: 	div_val = 32'h000002e8;
			45: 	div_val = 32'h000002d8;
			46: 	div_val = 32'h000002c8;
			47: 	div_val = 32'h000002b9;
			48: 	div_val = 32'h000002aa;
			49: 	div_val = 32'h0000029c;
			50: 	div_val = 32'h0000028f;
			51: 	div_val = 32'h00000282;
			52: 	div_val = 32'h00000276;
			53: 	div_val = 32'h0000026a;
			54: 	div_val = 32'h0000025e;
			55: 	div_val = 32'h00000253;
			56: 	div_val = 32'h00000249;
			57: 	div_val = 32'h0000023e;
			58: 	div_val = 32'h00000234;
			59: 	div_val = 32'h0000022b;
			60: 	div_val = 32'h00000222;
			61: 	div_val = 32'h00000219;
			62: 	div_val = 32'h00000210;
			63: 	div_val = 32'h00000208;
			64: 	div_val = 32'h00000200;
			65: 	div_val = 32'h000001f8;
			66: 	div_val = 32'h000001f0;
			67: 	div_val = 32'h000001e9;
			68: 	div_val = 32'h000001e1;
			69: 	div_val = 32'h000001da;
			70: 	div_val = 32'h000001d4;
			71: 	div_val = 32'h000001cd;
			72: 	div_val = 32'h000001c7;
			73: 	div_val = 32'h000001c0;
			74: 	div_val = 32'h000001ba;
			75: 	div_val = 32'h000001b4;
			76: 	div_val = 32'h000001af;
			77: 	div_val = 32'h000001a9;
			78: 	div_val = 32'h000001a4;
			79: 	div_val = 32'h0000019e;
			80: 	div_val = 32'h00000199;
			81: 	div_val = 32'h00000194;
			82: 	div_val = 32'h0000018f;
			83: 	div_val = 32'h0000018a;
			84: 	div_val = 32'h00000186;
			85: 	div_val = 32'h00000181;
			86: 	div_val = 32'h0000017d;
			87: 	div_val = 32'h00000178;
			88: 	div_val = 32'h00000174;
			89: 	div_val = 32'h00000170;
			90: 	div_val = 32'h0000016c;
			91: 	div_val = 32'h00000168;
			92: 	div_val = 32'h00000164;
			93: 	div_val = 32'h00000160;
			94: 	div_val = 32'h0000015c;
			95: 	div_val = 32'h00000158;
			96: 	div_val = 32'h00000155;
			97: 	div_val = 32'h00000151;
			98: 	div_val = 32'h0000014e;
			99: 	div_val = 32'h0000014a;
			100: 	div_val = 32'h00000147;
			101: 	div_val = 32'h00000144;
			102: 	div_val = 32'h00000141;
			103: 	div_val = 32'h0000013e;
			104: 	div_val = 32'h0000013b;
			105: 	div_val = 32'h00000138;
			106: 	div_val = 32'h00000135;
			107: 	div_val = 32'h00000132;
			108: 	div_val = 32'h0000012f;
			109: 	div_val = 32'h0000012c;
			110: 	div_val = 32'h00000129;
			111: 	div_val = 32'h00000127;
			112: 	div_val = 32'h00000124;
			113: 	div_val = 32'h00000121;
			114: 	div_val = 32'h0000011f;
			115: 	div_val = 32'h0000011c;
			116: 	div_val = 32'h0000011a;
			117: 	div_val = 32'h00000118;
			118: 	div_val = 32'h00000115;
			119: 	div_val = 32'h00000113;
			120: 	div_val = 32'h00000111;
			121: 	div_val = 32'h0000010e;
			122: 	div_val = 32'h0000010c;
			123: 	div_val = 32'h0000010a;
			124: 	div_val = 32'h00000108;
			125: 	div_val = 32'h00000106;
			126: 	div_val = 32'h00000104;
			127: 	div_val = 32'h00000102;
			default: div_val = 32'b0;
		endcase
	end
endmodule

module lut_256_divider
(	
	input logic [8:0] lut_sel,
	output logic signed[31:0] div_val
);
	always @(*) begin
		case(lut_sel)
			0: 	div_val = 32'b0;
			1: 	div_val = 32'd1 << 16;
			2: 	div_val = 32'h00004000;
			3: 	div_val = 32'h00002aaa;
			4: 	div_val = 32'h00002000;
			5: 	div_val = 32'h00001999;
			6: 	div_val = 32'h00001555;
			7: 	div_val = 32'h00001249;
			8: 	div_val = 32'h00001000;
			9: 	div_val = 32'h00000e38;
			10: 	div_val = 32'h00000ccc;
			11: 	div_val = 32'h00000ba2;
			12: 	div_val = 32'h00000aaa;
			13: 	div_val = 32'h000009d8;
			14: 	div_val = 32'h00000924;
			15: 	div_val = 32'h00000888;
			16: 	div_val = 32'h00000800;
			17: 	div_val = 32'h00000787;
			18: 	div_val = 32'h0000071c;
			19: 	div_val = 32'h000006bc;
			20: 	div_val = 32'h00000666;
			21: 	div_val = 32'h00000618;
			22: 	div_val = 32'h000005d1;
			23: 	div_val = 32'h00000590;
			24: 	div_val = 32'h00000555;
			25: 	div_val = 32'h0000051e;
			26: 	div_val = 32'h000004ec;
			27: 	div_val = 32'h000004bd;
			28: 	div_val = 32'h00000492;
			29: 	div_val = 32'h00000469;
			30: 	div_val = 32'h00000444;
			31: 	div_val = 32'h00000421;
			32: 	div_val = 32'h00000400;
			33: 	div_val = 32'h000003e0;
			34: 	div_val = 32'h000003c3;
			35: 	div_val = 32'h000003a8;
			36: 	div_val = 32'h0000038e;
			37: 	div_val = 32'h00000375;
			38: 	div_val = 32'h0000035e;
			39: 	div_val = 32'h00000348;
			40: 	div_val = 32'h00000333;
			41: 	div_val = 32'h0000031f;
			42: 	div_val = 32'h0000030c;
			43: 	div_val = 32'h000002fa;
			44: 	div_val = 32'h000002e8;
			45: 	div_val = 32'h000002d8;
			46: 	div_val = 32'h000002c8;
			47: 	div_val = 32'h000002b9;
			48: 	div_val = 32'h000002aa;
			49: 	div_val = 32'h0000029c;
			50: 	div_val = 32'h0000028f;
			51: 	div_val = 32'h00000282;
			52: 	div_val = 32'h00000276;
			53: 	div_val = 32'h0000026a;
			54: 	div_val = 32'h0000025e;
			55: 	div_val = 32'h00000253;
			56: 	div_val = 32'h00000249;
			57: 	div_val = 32'h0000023e;
			58: 	div_val = 32'h00000234;
			59: 	div_val = 32'h0000022b;
			60: 	div_val = 32'h00000222;
			61: 	div_val = 32'h00000219;
			62: 	div_val = 32'h00000210;
			63: 	div_val = 32'h00000208;
			64: 	div_val = 32'h00000200;
			65: 	div_val = 32'h000001f8;
			66: 	div_val = 32'h000001f0;
			67: 	div_val = 32'h000001e9;
			68: 	div_val = 32'h000001e1;
			69: 	div_val = 32'h000001da;
			70: 	div_val = 32'h000001d4;
			71: 	div_val = 32'h000001cd;
			72: 	div_val = 32'h000001c7;
			73: 	div_val = 32'h000001c0;
			74: 	div_val = 32'h000001ba;
			75: 	div_val = 32'h000001b4;
			76: 	div_val = 32'h000001af;
			77: 	div_val = 32'h000001a9;
			78: 	div_val = 32'h000001a4;
			79: 	div_val = 32'h0000019e;
			80: 	div_val = 32'h00000199;
			81: 	div_val = 32'h00000194;
			82: 	div_val = 32'h0000018f;
			83: 	div_val = 32'h0000018a;
			84: 	div_val = 32'h00000186;
			85: 	div_val = 32'h00000181;
			86: 	div_val = 32'h0000017d;
			87: 	div_val = 32'h00000178;
			88: 	div_val = 32'h00000174;
			89: 	div_val = 32'h00000170;
			90: 	div_val = 32'h0000016c;
			91: 	div_val = 32'h00000168;
			92: 	div_val = 32'h00000164;
			93: 	div_val = 32'h00000160;
			94: 	div_val = 32'h0000015c;
			95: 	div_val = 32'h00000158;
			96: 	div_val = 32'h00000155;
			97: 	div_val = 32'h00000151;
			98: 	div_val = 32'h0000014e;
			99: 	div_val = 32'h0000014a;
			100: 	div_val = 32'h00000147;
			101: 	div_val = 32'h00000144;
			102: 	div_val = 32'h00000141;
			103: 	div_val = 32'h0000013e;
			104: 	div_val = 32'h0000013b;
			105: 	div_val = 32'h00000138;
			106: 	div_val = 32'h00000135;
			107: 	div_val = 32'h00000132;
			108: 	div_val = 32'h0000012f;
			109: 	div_val = 32'h0000012c;
			110: 	div_val = 32'h00000129;
			111: 	div_val = 32'h00000127;
			112: 	div_val = 32'h00000124;
			113: 	div_val = 32'h00000121;
			114: 	div_val = 32'h0000011f;
			115: 	div_val = 32'h0000011c;
			116: 	div_val = 32'h0000011a;
			117: 	div_val = 32'h00000118;
			118: 	div_val = 32'h00000115;
			119: 	div_val = 32'h00000113;
			120: 	div_val = 32'h00000111;
			121: 	div_val = 32'h0000010e;
			122: 	div_val = 32'h0000010c;
			123: 	div_val = 32'h0000010a;
			124: 	div_val = 32'h00000108;
			125: 	div_val = 32'h00000106;
			126: 	div_val = 32'h00000104;
			127: 	div_val = 32'h00000102;
			128: 	div_val = 32'h00000100;
			129: 	div_val = 32'h000000fe;
			130: 	div_val = 32'h000000fc;
			131: 	div_val = 32'h000000fa;
			132: 	div_val = 32'h000000f8;
			133: 	div_val = 32'h000000f6;
			134: 	div_val = 32'h000000f4;
			135: 	div_val = 32'h000000f2;
			136: 	div_val = 32'h000000f0;
			137: 	div_val = 32'h000000ef;
			138: 	div_val = 32'h000000ed;
			139: 	div_val = 32'h000000eb;
			140: 	div_val = 32'h000000ea;
			141: 	div_val = 32'h000000e8;
			142: 	div_val = 32'h000000e6;
			143: 	div_val = 32'h000000e5;
			144: 	div_val = 32'h000000e3;
			145: 	div_val = 32'h000000e1;
			146: 	div_val = 32'h000000e0;
			147: 	div_val = 32'h000000de;
			148: 	div_val = 32'h000000dd;
			149: 	div_val = 32'h000000db;
			150: 	div_val = 32'h000000da;
			151: 	div_val = 32'h000000d9;
			152: 	div_val = 32'h000000d7;
			153: 	div_val = 32'h000000d6;
			154: 	div_val = 32'h000000d4;
			155: 	div_val = 32'h000000d3;
			156: 	div_val = 32'h000000d2;
			157: 	div_val = 32'h000000d0;
			158: 	div_val = 32'h000000cf;
			159: 	div_val = 32'h000000ce;
			160: 	div_val = 32'h000000cc;
			161: 	div_val = 32'h000000cb;
			162: 	div_val = 32'h000000ca;
			163: 	div_val = 32'h000000c9;
			164: 	div_val = 32'h000000c7;
			165: 	div_val = 32'h000000c6;
			166: 	div_val = 32'h000000c5;
			167: 	div_val = 32'h000000c4;
			168: 	div_val = 32'h000000c3;
			169: 	div_val = 32'h000000c1;
			170: 	div_val = 32'h000000c0;
			171: 	div_val = 32'h000000bf;
			172: 	div_val = 32'h000000be;
			173: 	div_val = 32'h000000bd;
			174: 	div_val = 32'h000000bc;
			175: 	div_val = 32'h000000bb;
			176: 	div_val = 32'h000000ba;
			177: 	div_val = 32'h000000b9;
			178: 	div_val = 32'h000000b8;
			179: 	div_val = 32'h000000b7;
			180: 	div_val = 32'h000000b6;
			181: 	div_val = 32'h000000b5;
			182: 	div_val = 32'h000000b4;
			183: 	div_val = 32'h000000b3;
			184: 	div_val = 32'h000000b2;
			185: 	div_val = 32'h000000b1;
			186: 	div_val = 32'h000000b0;
			187: 	div_val = 32'h000000af;
			188: 	div_val = 32'h000000ae;
			189: 	div_val = 32'h000000ad;
			190: 	div_val = 32'h000000ac;
			191: 	div_val = 32'h000000ab;
			192: 	div_val = 32'h000000aa;
			193: 	div_val = 32'h000000a9;
			194: 	div_val = 32'h000000a8;
			195: 	div_val = 32'h000000a8;
			196: 	div_val = 32'h000000a7;
			197: 	div_val = 32'h000000a6;
			198: 	div_val = 32'h000000a5;
			199: 	div_val = 32'h000000a4;
			200: 	div_val = 32'h000000a3;
			201: 	div_val = 32'h000000a3;
			202: 	div_val = 32'h000000a2;
			203: 	div_val = 32'h000000a1;
			204: 	div_val = 32'h000000a0;
			205: 	div_val = 32'h0000009f;
			206: 	div_val = 32'h0000009f;
			207: 	div_val = 32'h0000009e;
			208: 	div_val = 32'h0000009d;
			209: 	div_val = 32'h0000009c;
			210: 	div_val = 32'h0000009c;
			211: 	div_val = 32'h0000009b;
			212: 	div_val = 32'h0000009a;
			213: 	div_val = 32'h00000099;
			214: 	div_val = 32'h00000099;
			215: 	div_val = 32'h00000098;
			216: 	div_val = 32'h00000097;
			217: 	div_val = 32'h00000097;
			218: 	div_val = 32'h00000096;
			219: 	div_val = 32'h00000095;
			220: 	div_val = 32'h00000094;
			221: 	div_val = 32'h00000094;
			222: 	div_val = 32'h00000093;
			223: 	div_val = 32'h00000092;
			224: 	div_val = 32'h00000092;
			225: 	div_val = 32'h00000091;
			226: 	div_val = 32'h00000090;
			227: 	div_val = 32'h00000090;
			228: 	div_val = 32'h0000008f;
			229: 	div_val = 32'h0000008f;
			230: 	div_val = 32'h0000008e;
			231: 	div_val = 32'h0000008d;
			232: 	div_val = 32'h0000008d;
			233: 	div_val = 32'h0000008c;
			234: 	div_val = 32'h0000008c;
			235: 	div_val = 32'h0000008b;
			236: 	div_val = 32'h0000008a;
			237: 	div_val = 32'h0000008a;
			238: 	div_val = 32'h00000089;
			239: 	div_val = 32'h00000089;
			240: 	div_val = 32'h00000088;
			241: 	div_val = 32'h00000087;
			242: 	div_val = 32'h00000087;
			243: 	div_val = 32'h00000086;
			244: 	div_val = 32'h00000086;
			245: 	div_val = 32'h00000085;
			246: 	div_val = 32'h00000085;
			247: 	div_val = 32'h00000084;
			248: 	div_val = 32'h00000084;
			249: 	div_val = 32'h00000083;
			250: 	div_val = 32'h00000083;
			251: 	div_val = 32'h00000082;
			252: 	div_val = 32'h00000082;
			253: 	div_val = 32'h00000081;
			254: 	div_val = 32'h00000081;
			255: 	div_val = 32'h00000080;
			default: div_val = 32'b0;
		endcase
	end
endmodule

module lut_512_divider
(	
	input logic [9:0] lut_sel,
	output logic signed[31:0] div_val
);
	// Lookup table for values of lut_sel mapping to 1/lut_sel for values
	// from 1 to 31, and returning 0 for lut_sel = 0. This will lead to
	// the centering and matching factors being zeroed out if no neighboring boids are detected.
	
	always @(*) begin
		case(lut_sel)
			0: 	div_val = 32'b0;
			1: 	div_val = 32'd1 << 16;
			2: 	div_val = 32'h00004000;
			3: 	div_val = 32'h00002aaa;
			4: 	div_val = 32'h00002000;
			5: 	div_val = 32'h00001999;
			6: 	div_val = 32'h00001555;
			7: 	div_val = 32'h00001249;
			8: 	div_val = 32'h00001000;
			9: 	div_val = 32'h00000e38;
			10: 	div_val = 32'h00000ccc;
			11: 	div_val = 32'h00000ba2;
			12: 	div_val = 32'h00000aaa;
			13: 	div_val = 32'h000009d8;
			14: 	div_val = 32'h00000924;
			15: 	div_val = 32'h00000888;
			16: 	div_val = 32'h00000800;
			17: 	div_val = 32'h00000787;
			18: 	div_val = 32'h0000071c;
			19: 	div_val = 32'h000006bc;
			20: 	div_val = 32'h00000666;
			21: 	div_val = 32'h00000618;
			22: 	div_val = 32'h000005d1;
			23: 	div_val = 32'h00000590;
			24: 	div_val = 32'h00000555;
			25: 	div_val = 32'h0000051e;
			26: 	div_val = 32'h000004ec;
			27: 	div_val = 32'h000004bd;
			28: 	div_val = 32'h00000492;
			29: 	div_val = 32'h00000469;
			30: 	div_val = 32'h00000444;
			31: 	div_val = 32'h00000421;
			32: 	div_val = 32'h00000400;
			33: 	div_val = 32'h000003e0;
			34: 	div_val = 32'h000003c3;
			35: 	div_val = 32'h000003a8;
			36: 	div_val = 32'h0000038e;
			37: 	div_val = 32'h00000375;
			38: 	div_val = 32'h0000035e;
			39: 	div_val = 32'h00000348;
			40: 	div_val = 32'h00000333;
			41: 	div_val = 32'h0000031f;
			42: 	div_val = 32'h0000030c;
			43: 	div_val = 32'h000002fa;
			44: 	div_val = 32'h000002e8;
			45: 	div_val = 32'h000002d8;
			46: 	div_val = 32'h000002c8;
			47: 	div_val = 32'h000002b9;
			48: 	div_val = 32'h000002aa;
			49: 	div_val = 32'h0000029c;
			50: 	div_val = 32'h0000028f;
			51: 	div_val = 32'h00000282;
			52: 	div_val = 32'h00000276;
			53: 	div_val = 32'h0000026a;
			54: 	div_val = 32'h0000025e;
			55: 	div_val = 32'h00000253;
			56: 	div_val = 32'h00000249;
			57: 	div_val = 32'h0000023e;
			58: 	div_val = 32'h00000234;
			59: 	div_val = 32'h0000022b;
			60: 	div_val = 32'h00000222;
			61: 	div_val = 32'h00000219;
			62: 	div_val = 32'h00000210;
			63: 	div_val = 32'h00000208;
			64: 	div_val = 32'h00000200;
			65: 	div_val = 32'h000001f8;
			66: 	div_val = 32'h000001f0;
			67: 	div_val = 32'h000001e9;
			68: 	div_val = 32'h000001e1;
			69: 	div_val = 32'h000001da;
			70: 	div_val = 32'h000001d4;
			71: 	div_val = 32'h000001cd;
			72: 	div_val = 32'h000001c7;
			73: 	div_val = 32'h000001c0;
			74: 	div_val = 32'h000001ba;
			75: 	div_val = 32'h000001b4;
			76: 	div_val = 32'h000001af;
			77: 	div_val = 32'h000001a9;
			78: 	div_val = 32'h000001a4;
			79: 	div_val = 32'h0000019e;
			80: 	div_val = 32'h00000199;
			81: 	div_val = 32'h00000194;
			82: 	div_val = 32'h0000018f;
			83: 	div_val = 32'h0000018a;
			84: 	div_val = 32'h00000186;
			85: 	div_val = 32'h00000181;
			86: 	div_val = 32'h0000017d;
			87: 	div_val = 32'h00000178;
			88: 	div_val = 32'h00000174;
			89: 	div_val = 32'h00000170;
			90: 	div_val = 32'h0000016c;
			91: 	div_val = 32'h00000168;
			92: 	div_val = 32'h00000164;
			93: 	div_val = 32'h00000160;
			94: 	div_val = 32'h0000015c;
			95: 	div_val = 32'h00000158;
			96: 	div_val = 32'h00000155;
			97: 	div_val = 32'h00000151;
			98: 	div_val = 32'h0000014e;
			99: 	div_val = 32'h0000014a;
			100: 	div_val = 32'h00000147;
			101: 	div_val = 32'h00000144;
			102: 	div_val = 32'h00000141;
			103: 	div_val = 32'h0000013e;
			104: 	div_val = 32'h0000013b;
			105: 	div_val = 32'h00000138;
			106: 	div_val = 32'h00000135;
			107: 	div_val = 32'h00000132;
			108: 	div_val = 32'h0000012f;
			109: 	div_val = 32'h0000012c;
			110: 	div_val = 32'h00000129;
			111: 	div_val = 32'h00000127;
			112: 	div_val = 32'h00000124;
			113: 	div_val = 32'h00000121;
			114: 	div_val = 32'h0000011f;
			115: 	div_val = 32'h0000011c;
			116: 	div_val = 32'h0000011a;
			117: 	div_val = 32'h00000118;
			118: 	div_val = 32'h00000115;
			119: 	div_val = 32'h00000113;
			120: 	div_val = 32'h00000111;
			121: 	div_val = 32'h0000010e;
			122: 	div_val = 32'h0000010c;
			123: 	div_val = 32'h0000010a;
			124: 	div_val = 32'h00000108;
			125: 	div_val = 32'h00000106;
			126: 	div_val = 32'h00000104;
			127: 	div_val = 32'h00000102;
			128: 	div_val = 32'h00000100;
			129: 	div_val = 32'h000000fe;
			130: 	div_val = 32'h000000fc;
			131: 	div_val = 32'h000000fa;
			132: 	div_val = 32'h000000f8;
			133: 	div_val = 32'h000000f6;
			134: 	div_val = 32'h000000f4;
			135: 	div_val = 32'h000000f2;
			136: 	div_val = 32'h000000f0;
			137: 	div_val = 32'h000000ef;
			138: 	div_val = 32'h000000ed;
			139: 	div_val = 32'h000000eb;
			140: 	div_val = 32'h000000ea;
			141: 	div_val = 32'h000000e8;
			142: 	div_val = 32'h000000e6;
			143: 	div_val = 32'h000000e5;
			144: 	div_val = 32'h000000e3;
			145: 	div_val = 32'h000000e1;
			146: 	div_val = 32'h000000e0;
			147: 	div_val = 32'h000000de;
			148: 	div_val = 32'h000000dd;
			149: 	div_val = 32'h000000db;
			150: 	div_val = 32'h000000da;
			151: 	div_val = 32'h000000d9;
			152: 	div_val = 32'h000000d7;
			153: 	div_val = 32'h000000d6;
			154: 	div_val = 32'h000000d4;
			155: 	div_val = 32'h000000d3;
			156: 	div_val = 32'h000000d2;
			157: 	div_val = 32'h000000d0;
			158: 	div_val = 32'h000000cf;
			159: 	div_val = 32'h000000ce;
			160: 	div_val = 32'h000000cc;
			161: 	div_val = 32'h000000cb;
			162: 	div_val = 32'h000000ca;
			163: 	div_val = 32'h000000c9;
			164: 	div_val = 32'h000000c7;
			165: 	div_val = 32'h000000c6;
			166: 	div_val = 32'h000000c5;
			167: 	div_val = 32'h000000c4;
			168: 	div_val = 32'h000000c3;
			169: 	div_val = 32'h000000c1;
			170: 	div_val = 32'h000000c0;
			171: 	div_val = 32'h000000bf;
			172: 	div_val = 32'h000000be;
			173: 	div_val = 32'h000000bd;
			174: 	div_val = 32'h000000bc;
			175: 	div_val = 32'h000000bb;
			176: 	div_val = 32'h000000ba;
			177: 	div_val = 32'h000000b9;
			178: 	div_val = 32'h000000b8;
			179: 	div_val = 32'h000000b7;
			180: 	div_val = 32'h000000b6;
			181: 	div_val = 32'h000000b5;
			182: 	div_val = 32'h000000b4;
			183: 	div_val = 32'h000000b3;
			184: 	div_val = 32'h000000b2;
			185: 	div_val = 32'h000000b1;
			186: 	div_val = 32'h000000b0;
			187: 	div_val = 32'h000000af;
			188: 	div_val = 32'h000000ae;
			189: 	div_val = 32'h000000ad;
			190: 	div_val = 32'h000000ac;
			191: 	div_val = 32'h000000ab;
			192: 	div_val = 32'h000000aa;
			193: 	div_val = 32'h000000a9;
			194: 	div_val = 32'h000000a8;
			195: 	div_val = 32'h000000a8;
			196: 	div_val = 32'h000000a7;
			197: 	div_val = 32'h000000a6;
			198: 	div_val = 32'h000000a5;
			199: 	div_val = 32'h000000a4;
			200: 	div_val = 32'h000000a3;
			201: 	div_val = 32'h000000a3;
			202: 	div_val = 32'h000000a2;
			203: 	div_val = 32'h000000a1;
			204: 	div_val = 32'h000000a0;
			205: 	div_val = 32'h0000009f;
			206: 	div_val = 32'h0000009f;
			207: 	div_val = 32'h0000009e;
			208: 	div_val = 32'h0000009d;
			209: 	div_val = 32'h0000009c;
			210: 	div_val = 32'h0000009c;
			211: 	div_val = 32'h0000009b;
			212: 	div_val = 32'h0000009a;
			213: 	div_val = 32'h00000099;
			214: 	div_val = 32'h00000099;
			215: 	div_val = 32'h00000098;
			216: 	div_val = 32'h00000097;
			217: 	div_val = 32'h00000097;
			218: 	div_val = 32'h00000096;
			219: 	div_val = 32'h00000095;
			220: 	div_val = 32'h00000094;
			221: 	div_val = 32'h00000094;
			222: 	div_val = 32'h00000093;
			223: 	div_val = 32'h00000092;
			224: 	div_val = 32'h00000092;
			225: 	div_val = 32'h00000091;
			226: 	div_val = 32'h00000090;
			227: 	div_val = 32'h00000090;
			228: 	div_val = 32'h0000008f;
			229: 	div_val = 32'h0000008f;
			230: 	div_val = 32'h0000008e;
			231: 	div_val = 32'h0000008d;
			232: 	div_val = 32'h0000008d;
			233: 	div_val = 32'h0000008c;
			234: 	div_val = 32'h0000008c;
			235: 	div_val = 32'h0000008b;
			236: 	div_val = 32'h0000008a;
			237: 	div_val = 32'h0000008a;
			238: 	div_val = 32'h00000089;
			239: 	div_val = 32'h00000089;
			240: 	div_val = 32'h00000088;
			241: 	div_val = 32'h00000087;
			242: 	div_val = 32'h00000087;
			243: 	div_val = 32'h00000086;
			244: 	div_val = 32'h00000086;
			245: 	div_val = 32'h00000085;
			246: 	div_val = 32'h00000085;
			247: 	div_val = 32'h00000084;
			248: 	div_val = 32'h00000084;
			249: 	div_val = 32'h00000083;
			250: 	div_val = 32'h00000083;
			251: 	div_val = 32'h00000082;
			252: 	div_val = 32'h00000082;
			253: 	div_val = 32'h00000081;
			254: 	div_val = 32'h00000081;
			255: 	div_val = 32'h00000080;
			256: 	div_val = 32'h00000080;
			257: 	div_val = 32'h0000007f;
			258: 	div_val = 32'h0000007f;
			259: 	div_val = 32'h0000007e;
			260: 	div_val = 32'h0000007e;
			261: 	div_val = 32'h0000007d;
			262: 	div_val = 32'h0000007d;
			263: 	div_val = 32'h0000007c;
			264: 	div_val = 32'h0000007c;
			265: 	div_val = 32'h0000007b;
			266: 	div_val = 32'h0000007b;
			267: 	div_val = 32'h0000007a;
			268: 	div_val = 32'h0000007a;
			269: 	div_val = 32'h00000079;
			270: 	div_val = 32'h00000079;
			271: 	div_val = 32'h00000078;
			272: 	div_val = 32'h00000078;
			273: 	div_val = 32'h00000078;
			274: 	div_val = 32'h00000077;
			275: 	div_val = 32'h00000077;
			276: 	div_val = 32'h00000076;
			277: 	div_val = 32'h00000076;
			278: 	div_val = 32'h00000075;
			279: 	div_val = 32'h00000075;
			280: 	div_val = 32'h00000075;
			281: 	div_val = 32'h00000074;
			282: 	div_val = 32'h00000074;
			283: 	div_val = 32'h00000073;
			284: 	div_val = 32'h00000073;
			285: 	div_val = 32'h00000072;
			286: 	div_val = 32'h00000072;
			287: 	div_val = 32'h00000072;
			288: 	div_val = 32'h00000071;
			289: 	div_val = 32'h00000071;
			290: 	div_val = 32'h00000070;
			291: 	div_val = 32'h00000070;
			292: 	div_val = 32'h00000070;
			293: 	div_val = 32'h0000006f;
			294: 	div_val = 32'h0000006f;
			295: 	div_val = 32'h0000006f;
			296: 	div_val = 32'h0000006e;
			297: 	div_val = 32'h0000006e;
			298: 	div_val = 32'h0000006d;
			299: 	div_val = 32'h0000006d;
			300: 	div_val = 32'h0000006d;
			301: 	div_val = 32'h0000006c;
			302: 	div_val = 32'h0000006c;
			303: 	div_val = 32'h0000006c;
			304: 	div_val = 32'h0000006b;
			305: 	div_val = 32'h0000006b;
			306: 	div_val = 32'h0000006b;
			307: 	div_val = 32'h0000006a;
			308: 	div_val = 32'h0000006a;
			309: 	div_val = 32'h0000006a;
			310: 	div_val = 32'h00000069;
			311: 	div_val = 32'h00000069;
			312: 	div_val = 32'h00000069;
			313: 	div_val = 32'h00000068;
			314: 	div_val = 32'h00000068;
			315: 	div_val = 32'h00000068;
			316: 	div_val = 32'h00000067;
			317: 	div_val = 32'h00000067;
			318: 	div_val = 32'h00000067;
			319: 	div_val = 32'h00000066;
			320: 	div_val = 32'h00000066;
			321: 	div_val = 32'h00000066;
			322: 	div_val = 32'h00000065;
			323: 	div_val = 32'h00000065;
			324: 	div_val = 32'h00000065;
			325: 	div_val = 32'h00000064;
			326: 	div_val = 32'h00000064;
			327: 	div_val = 32'h00000064;
			328: 	div_val = 32'h00000063;
			329: 	div_val = 32'h00000063;
			330: 	div_val = 32'h00000063;
			331: 	div_val = 32'h00000062;
			332: 	div_val = 32'h00000062;
			333: 	div_val = 32'h00000062;
			334: 	div_val = 32'h00000062;
			335: 	div_val = 32'h00000061;
			336: 	div_val = 32'h00000061;
			337: 	div_val = 32'h00000061;
			338: 	div_val = 32'h00000060;
			339: 	div_val = 32'h00000060;
			340: 	div_val = 32'h00000060;
			341: 	div_val = 32'h00000060;
			342: 	div_val = 32'h0000005f;
			343: 	div_val = 32'h0000005f;
			344: 	div_val = 32'h0000005f;
			345: 	div_val = 32'h0000005e;
			346: 	div_val = 32'h0000005e;
			347: 	div_val = 32'h0000005e;
			348: 	div_val = 32'h0000005e;
			349: 	div_val = 32'h0000005d;
			350: 	div_val = 32'h0000005d;
			351: 	div_val = 32'h0000005d;
			352: 	div_val = 32'h0000005d;
			353: 	div_val = 32'h0000005c;
			354: 	div_val = 32'h0000005c;
			355: 	div_val = 32'h0000005c;
			356: 	div_val = 32'h0000005c;
			357: 	div_val = 32'h0000005b;
			358: 	div_val = 32'h0000005b;
			359: 	div_val = 32'h0000005b;
			360: 	div_val = 32'h0000005b;
			361: 	div_val = 32'h0000005a;
			362: 	div_val = 32'h0000005a;
			363: 	div_val = 32'h0000005a;
			364: 	div_val = 32'h0000005a;
			365: 	div_val = 32'h00000059;
			366: 	div_val = 32'h00000059;
			367: 	div_val = 32'h00000059;
			368: 	div_val = 32'h00000059;
			369: 	div_val = 32'h00000058;
			370: 	div_val = 32'h00000058;
			371: 	div_val = 32'h00000058;
			372: 	div_val = 32'h00000058;
			373: 	div_val = 32'h00000057;
			374: 	div_val = 32'h00000057;
			375: 	div_val = 32'h00000057;
			376: 	div_val = 32'h00000057;
			377: 	div_val = 32'h00000056;
			378: 	div_val = 32'h00000056;
			379: 	div_val = 32'h00000056;
			380: 	div_val = 32'h00000056;
			381: 	div_val = 32'h00000056;
			382: 	div_val = 32'h00000055;
			383: 	div_val = 32'h00000055;
			384: 	div_val = 32'h00000055;
			385: 	div_val = 32'h00000055;
			386: 	div_val = 32'h00000054;
			387: 	div_val = 32'h00000054;
			388: 	div_val = 32'h00000054;
			389: 	div_val = 32'h00000054;
			390: 	div_val = 32'h00000054;
			391: 	div_val = 32'h00000053;
			392: 	div_val = 32'h00000053;
			393: 	div_val = 32'h00000053;
			394: 	div_val = 32'h00000053;
			395: 	div_val = 32'h00000052;
			396: 	div_val = 32'h00000052;
			397: 	div_val = 32'h00000052;
			398: 	div_val = 32'h00000052;
			399: 	div_val = 32'h00000052;
			400: 	div_val = 32'h00000051;
			401: 	div_val = 32'h00000051;
			402: 	div_val = 32'h00000051;
			403: 	div_val = 32'h00000051;
			404: 	div_val = 32'h00000051;
			405: 	div_val = 32'h00000050;
			406: 	div_val = 32'h00000050;
			407: 	div_val = 32'h00000050;
			408: 	div_val = 32'h00000050;
			409: 	div_val = 32'h00000050;
			410: 	div_val = 32'h0000004f;
			411: 	div_val = 32'h0000004f;
			412: 	div_val = 32'h0000004f;
			413: 	div_val = 32'h0000004f;
			414: 	div_val = 32'h0000004f;
			415: 	div_val = 32'h0000004e;
			416: 	div_val = 32'h0000004e;
			417: 	div_val = 32'h0000004e;
			418: 	div_val = 32'h0000004e;
			419: 	div_val = 32'h0000004e;
			420: 	div_val = 32'h0000004e;
			421: 	div_val = 32'h0000004d;
			422: 	div_val = 32'h0000004d;
			423: 	div_val = 32'h0000004d;
			424: 	div_val = 32'h0000004d;
			425: 	div_val = 32'h0000004d;
			426: 	div_val = 32'h0000004c;
			427: 	div_val = 32'h0000004c;
			428: 	div_val = 32'h0000004c;
			429: 	div_val = 32'h0000004c;
			430: 	div_val = 32'h0000004c;
			431: 	div_val = 32'h0000004c;
			432: 	div_val = 32'h0000004b;
			433: 	div_val = 32'h0000004b;
			434: 	div_val = 32'h0000004b;
			435: 	div_val = 32'h0000004b;
			436: 	div_val = 32'h0000004b;
			437: 	div_val = 32'h0000004a;
			438: 	div_val = 32'h0000004a;
			439: 	div_val = 32'h0000004a;
			440: 	div_val = 32'h0000004a;
			441: 	div_val = 32'h0000004a;
			442: 	div_val = 32'h0000004a;
			443: 	div_val = 32'h00000049;
			444: 	div_val = 32'h00000049;
			445: 	div_val = 32'h00000049;
			446: 	div_val = 32'h00000049;
			447: 	div_val = 32'h00000049;
			448: 	div_val = 32'h00000049;
			449: 	div_val = 32'h00000048;
			450: 	div_val = 32'h00000048;
			451: 	div_val = 32'h00000048;
			452: 	div_val = 32'h00000048;
			453: 	div_val = 32'h00000048;
			454: 	div_val = 32'h00000048;
			455: 	div_val = 32'h00000048;
			456: 	div_val = 32'h00000047;
			457: 	div_val = 32'h00000047;
			458: 	div_val = 32'h00000047;
			459: 	div_val = 32'h00000047;
			460: 	div_val = 32'h00000047;
			461: 	div_val = 32'h00000047;
			462: 	div_val = 32'h00000046;
			463: 	div_val = 32'h00000046;
			464: 	div_val = 32'h00000046;
			465: 	div_val = 32'h00000046;
			466: 	div_val = 32'h00000046;
			467: 	div_val = 32'h00000046;
			468: 	div_val = 32'h00000046;
			469: 	div_val = 32'h00000045;
			470: 	div_val = 32'h00000045;
			471: 	div_val = 32'h00000045;
			472: 	div_val = 32'h00000045;
			473: 	div_val = 32'h00000045;
			474: 	div_val = 32'h00000045;
			475: 	div_val = 32'h00000044;
			476: 	div_val = 32'h00000044;
			477: 	div_val = 32'h00000044;
			478: 	div_val = 32'h00000044;
			479: 	div_val = 32'h00000044;
			480: 	div_val = 32'h00000044;
			481: 	div_val = 32'h00000044;
			482: 	div_val = 32'h00000043;
			483: 	div_val = 32'h00000043;
			484: 	div_val = 32'h00000043;
			485: 	div_val = 32'h00000043;
			486: 	div_val = 32'h00000043;
			487: 	div_val = 32'h00000043;
			488: 	div_val = 32'h00000043;
			489: 	div_val = 32'h00000043;
			490: 	div_val = 32'h00000042;
			491: 	div_val = 32'h00000042;
			492: 	div_val = 32'h00000042;
			493: 	div_val = 32'h00000042;
			494: 	div_val = 32'h00000042;
			495: 	div_val = 32'h00000042;
			496: 	div_val = 32'h00000042;
			497: 	div_val = 32'h00000041;
			498: 	div_val = 32'h00000041;
			499: 	div_val = 32'h00000041;
			500: 	div_val = 32'h00000041;
			501: 	div_val = 32'h00000041;
			502: 	div_val = 32'h00000041;
			503: 	div_val = 32'h00000041;
			504: 	div_val = 32'h00000041;
			505: 	div_val = 32'h00000040;
			506: 	div_val = 32'h00000040;
			507: 	div_val = 32'h00000040;
			508: 	div_val = 32'h00000040;
			509: 	div_val = 32'h00000040;
			510: 	div_val = 32'h00000040;
			511: 	div_val = 32'h00000040;
			default: div_val = 32'b0;
		endcase
	end

endmodule

module lut_1024_divider
(	
	input logic [10:0] lut_sel,
	output logic signed[31:0] div_val
);
	// Lookup table for values of lut_sel mapping to 1/lut_sel for values
	// from 1 to 31, and returning 0 for lut_sel = 0. This will lead to
	// the centering and matching factors being zeroed out if no neighboring boids are detected.
	
	always @(*) begin
		case(lut_sel)
			0: 	div_val = 32'b0;
			1: 	div_val = 32'd1 << 16;
			2: 	div_val = 32'h00004000;
			3: 	div_val = 32'h00002aaa;
			4: 	div_val = 32'h00002000;
			5: 	div_val = 32'h00001999;
			6: 	div_val = 32'h00001555;
			7: 	div_val = 32'h00001249;
			8: 	div_val = 32'h00001000;
			9: 	div_val = 32'h00000e38;
			10: 	div_val = 32'h00000ccc;
			11: 	div_val = 32'h00000ba2;
			12: 	div_val = 32'h00000aaa;
			13: 	div_val = 32'h000009d8;
			14: 	div_val = 32'h00000924;
			15: 	div_val = 32'h00000888;
			16: 	div_val = 32'h00000800;
			17: 	div_val = 32'h00000787;
			18: 	div_val = 32'h0000071c;
			19: 	div_val = 32'h000006bc;
			20: 	div_val = 32'h00000666;
			21: 	div_val = 32'h00000618;
			22: 	div_val = 32'h000005d1;
			23: 	div_val = 32'h00000590;
			24: 	div_val = 32'h00000555;
			25: 	div_val = 32'h0000051e;
			26: 	div_val = 32'h000004ec;
			27: 	div_val = 32'h000004bd;
			28: 	div_val = 32'h00000492;
			29: 	div_val = 32'h00000469;
			30: 	div_val = 32'h00000444;
			31: 	div_val = 32'h00000421;
			32: 	div_val = 32'h00000400;
			33: 	div_val = 32'h000003e0;
			34: 	div_val = 32'h000003c3;
			35: 	div_val = 32'h000003a8;
			36: 	div_val = 32'h0000038e;
			37: 	div_val = 32'h00000375;
			38: 	div_val = 32'h0000035e;
			39: 	div_val = 32'h00000348;
			40: 	div_val = 32'h00000333;
			41: 	div_val = 32'h0000031f;
			42: 	div_val = 32'h0000030c;
			43: 	div_val = 32'h000002fa;
			44: 	div_val = 32'h000002e8;
			45: 	div_val = 32'h000002d8;
			46: 	div_val = 32'h000002c8;
			47: 	div_val = 32'h000002b9;
			48: 	div_val = 32'h000002aa;
			49: 	div_val = 32'h0000029c;
			50: 	div_val = 32'h0000028f;
			51: 	div_val = 32'h00000282;
			52: 	div_val = 32'h00000276;
			53: 	div_val = 32'h0000026a;
			54: 	div_val = 32'h0000025e;
			55: 	div_val = 32'h00000253;
			56: 	div_val = 32'h00000249;
			57: 	div_val = 32'h0000023e;
			58: 	div_val = 32'h00000234;
			59: 	div_val = 32'h0000022b;
			60: 	div_val = 32'h00000222;
			61: 	div_val = 32'h00000219;
			62: 	div_val = 32'h00000210;
			63: 	div_val = 32'h00000208;
			64: 	div_val = 32'h00000200;
			65: 	div_val = 32'h000001f8;
			66: 	div_val = 32'h000001f0;
			67: 	div_val = 32'h000001e9;
			68: 	div_val = 32'h000001e1;
			69: 	div_val = 32'h000001da;
			70: 	div_val = 32'h000001d4;
			71: 	div_val = 32'h000001cd;
			72: 	div_val = 32'h000001c7;
			73: 	div_val = 32'h000001c0;
			74: 	div_val = 32'h000001ba;
			75: 	div_val = 32'h000001b4;
			76: 	div_val = 32'h000001af;
			77: 	div_val = 32'h000001a9;
			78: 	div_val = 32'h000001a4;
			79: 	div_val = 32'h0000019e;
			80: 	div_val = 32'h00000199;
			81: 	div_val = 32'h00000194;
			82: 	div_val = 32'h0000018f;
			83: 	div_val = 32'h0000018a;
			84: 	div_val = 32'h00000186;
			85: 	div_val = 32'h00000181;
			86: 	div_val = 32'h0000017d;
			87: 	div_val = 32'h00000178;
			88: 	div_val = 32'h00000174;
			89: 	div_val = 32'h00000170;
			90: 	div_val = 32'h0000016c;
			91: 	div_val = 32'h00000168;
			92: 	div_val = 32'h00000164;
			93: 	div_val = 32'h00000160;
			94: 	div_val = 32'h0000015c;
			95: 	div_val = 32'h00000158;
			96: 	div_val = 32'h00000155;
			97: 	div_val = 32'h00000151;
			98: 	div_val = 32'h0000014e;
			99: 	div_val = 32'h0000014a;
			100: 	div_val = 32'h00000147;
			101: 	div_val = 32'h00000144;
			102: 	div_val = 32'h00000141;
			103: 	div_val = 32'h0000013e;
			104: 	div_val = 32'h0000013b;
			105: 	div_val = 32'h00000138;
			106: 	div_val = 32'h00000135;
			107: 	div_val = 32'h00000132;
			108: 	div_val = 32'h0000012f;
			109: 	div_val = 32'h0000012c;
			110: 	div_val = 32'h00000129;
			111: 	div_val = 32'h00000127;
			112: 	div_val = 32'h00000124;
			113: 	div_val = 32'h00000121;
			114: 	div_val = 32'h0000011f;
			115: 	div_val = 32'h0000011c;
			116: 	div_val = 32'h0000011a;
			117: 	div_val = 32'h00000118;
			118: 	div_val = 32'h00000115;
			119: 	div_val = 32'h00000113;
			120: 	div_val = 32'h00000111;
			121: 	div_val = 32'h0000010e;
			122: 	div_val = 32'h0000010c;
			123: 	div_val = 32'h0000010a;
			124: 	div_val = 32'h00000108;
			125: 	div_val = 32'h00000106;
			126: 	div_val = 32'h00000104;
			127: 	div_val = 32'h00000102;
			128: 	div_val = 32'h00000100;
			129: 	div_val = 32'h000000fe;
			130: 	div_val = 32'h000000fc;
			131: 	div_val = 32'h000000fa;
			132: 	div_val = 32'h000000f8;
			133: 	div_val = 32'h000000f6;
			134: 	div_val = 32'h000000f4;
			135: 	div_val = 32'h000000f2;
			136: 	div_val = 32'h000000f0;
			137: 	div_val = 32'h000000ef;
			138: 	div_val = 32'h000000ed;
			139: 	div_val = 32'h000000eb;
			140: 	div_val = 32'h000000ea;
			141: 	div_val = 32'h000000e8;
			142: 	div_val = 32'h000000e6;
			143: 	div_val = 32'h000000e5;
			144: 	div_val = 32'h000000e3;
			145: 	div_val = 32'h000000e1;
			146: 	div_val = 32'h000000e0;
			147: 	div_val = 32'h000000de;
			148: 	div_val = 32'h000000dd;
			149: 	div_val = 32'h000000db;
			150: 	div_val = 32'h000000da;
			151: 	div_val = 32'h000000d9;
			152: 	div_val = 32'h000000d7;
			153: 	div_val = 32'h000000d6;
			154: 	div_val = 32'h000000d4;
			155: 	div_val = 32'h000000d3;
			156: 	div_val = 32'h000000d2;
			157: 	div_val = 32'h000000d0;
			158: 	div_val = 32'h000000cf;
			159: 	div_val = 32'h000000ce;
			160: 	div_val = 32'h000000cc;
			161: 	div_val = 32'h000000cb;
			162: 	div_val = 32'h000000ca;
			163: 	div_val = 32'h000000c9;
			164: 	div_val = 32'h000000c7;
			165: 	div_val = 32'h000000c6;
			166: 	div_val = 32'h000000c5;
			167: 	div_val = 32'h000000c4;
			168: 	div_val = 32'h000000c3;
			169: 	div_val = 32'h000000c1;
			170: 	div_val = 32'h000000c0;
			171: 	div_val = 32'h000000bf;
			172: 	div_val = 32'h000000be;
			173: 	div_val = 32'h000000bd;
			174: 	div_val = 32'h000000bc;
			175: 	div_val = 32'h000000bb;
			176: 	div_val = 32'h000000ba;
			177: 	div_val = 32'h000000b9;
			178: 	div_val = 32'h000000b8;
			179: 	div_val = 32'h000000b7;
			180: 	div_val = 32'h000000b6;
			181: 	div_val = 32'h000000b5;
			182: 	div_val = 32'h000000b4;
			183: 	div_val = 32'h000000b3;
			184: 	div_val = 32'h000000b2;
			185: 	div_val = 32'h000000b1;
			186: 	div_val = 32'h000000b0;
			187: 	div_val = 32'h000000af;
			188: 	div_val = 32'h000000ae;
			189: 	div_val = 32'h000000ad;
			190: 	div_val = 32'h000000ac;
			191: 	div_val = 32'h000000ab;
			192: 	div_val = 32'h000000aa;
			193: 	div_val = 32'h000000a9;
			194: 	div_val = 32'h000000a8;
			195: 	div_val = 32'h000000a8;
			196: 	div_val = 32'h000000a7;
			197: 	div_val = 32'h000000a6;
			198: 	div_val = 32'h000000a5;
			199: 	div_val = 32'h000000a4;
			200: 	div_val = 32'h000000a3;
			201: 	div_val = 32'h000000a3;
			202: 	div_val = 32'h000000a2;
			203: 	div_val = 32'h000000a1;
			204: 	div_val = 32'h000000a0;
			205: 	div_val = 32'h0000009f;
			206: 	div_val = 32'h0000009f;
			207: 	div_val = 32'h0000009e;
			208: 	div_val = 32'h0000009d;
			209: 	div_val = 32'h0000009c;
			210: 	div_val = 32'h0000009c;
			211: 	div_val = 32'h0000009b;
			212: 	div_val = 32'h0000009a;
			213: 	div_val = 32'h00000099;
			214: 	div_val = 32'h00000099;
			215: 	div_val = 32'h00000098;
			216: 	div_val = 32'h00000097;
			217: 	div_val = 32'h00000097;
			218: 	div_val = 32'h00000096;
			219: 	div_val = 32'h00000095;
			220: 	div_val = 32'h00000094;
			221: 	div_val = 32'h00000094;
			222: 	div_val = 32'h00000093;
			223: 	div_val = 32'h00000092;
			224: 	div_val = 32'h00000092;
			225: 	div_val = 32'h00000091;
			226: 	div_val = 32'h00000090;
			227: 	div_val = 32'h00000090;
			228: 	div_val = 32'h0000008f;
			229: 	div_val = 32'h0000008f;
			230: 	div_val = 32'h0000008e;
			231: 	div_val = 32'h0000008d;
			232: 	div_val = 32'h0000008d;
			233: 	div_val = 32'h0000008c;
			234: 	div_val = 32'h0000008c;
			235: 	div_val = 32'h0000008b;
			236: 	div_val = 32'h0000008a;
			237: 	div_val = 32'h0000008a;
			238: 	div_val = 32'h00000089;
			239: 	div_val = 32'h00000089;
			240: 	div_val = 32'h00000088;
			241: 	div_val = 32'h00000087;
			242: 	div_val = 32'h00000087;
			243: 	div_val = 32'h00000086;
			244: 	div_val = 32'h00000086;
			245: 	div_val = 32'h00000085;
			246: 	div_val = 32'h00000085;
			247: 	div_val = 32'h00000084;
			248: 	div_val = 32'h00000084;
			249: 	div_val = 32'h00000083;
			250: 	div_val = 32'h00000083;
			251: 	div_val = 32'h00000082;
			252: 	div_val = 32'h00000082;
			253: 	div_val = 32'h00000081;
			254: 	div_val = 32'h00000081;
			255: 	div_val = 32'h00000080;
			256: 	div_val = 32'h00000080;
			257: 	div_val = 32'h0000007f;
			258: 	div_val = 32'h0000007f;
			259: 	div_val = 32'h0000007e;
			260: 	div_val = 32'h0000007e;
			261: 	div_val = 32'h0000007d;
			262: 	div_val = 32'h0000007d;
			263: 	div_val = 32'h0000007c;
			264: 	div_val = 32'h0000007c;
			265: 	div_val = 32'h0000007b;
			266: 	div_val = 32'h0000007b;
			267: 	div_val = 32'h0000007a;
			268: 	div_val = 32'h0000007a;
			269: 	div_val = 32'h00000079;
			270: 	div_val = 32'h00000079;
			271: 	div_val = 32'h00000078;
			272: 	div_val = 32'h00000078;
			273: 	div_val = 32'h00000078;
			274: 	div_val = 32'h00000077;
			275: 	div_val = 32'h00000077;
			276: 	div_val = 32'h00000076;
			277: 	div_val = 32'h00000076;
			278: 	div_val = 32'h00000075;
			279: 	div_val = 32'h00000075;
			280: 	div_val = 32'h00000075;
			281: 	div_val = 32'h00000074;
			282: 	div_val = 32'h00000074;
			283: 	div_val = 32'h00000073;
			284: 	div_val = 32'h00000073;
			285: 	div_val = 32'h00000072;
			286: 	div_val = 32'h00000072;
			287: 	div_val = 32'h00000072;
			288: 	div_val = 32'h00000071;
			289: 	div_val = 32'h00000071;
			290: 	div_val = 32'h00000070;
			291: 	div_val = 32'h00000070;
			292: 	div_val = 32'h00000070;
			293: 	div_val = 32'h0000006f;
			294: 	div_val = 32'h0000006f;
			295: 	div_val = 32'h0000006f;
			296: 	div_val = 32'h0000006e;
			297: 	div_val = 32'h0000006e;
			298: 	div_val = 32'h0000006d;
			299: 	div_val = 32'h0000006d;
			300: 	div_val = 32'h0000006d;
			301: 	div_val = 32'h0000006c;
			302: 	div_val = 32'h0000006c;
			303: 	div_val = 32'h0000006c;
			304: 	div_val = 32'h0000006b;
			305: 	div_val = 32'h0000006b;
			306: 	div_val = 32'h0000006b;
			307: 	div_val = 32'h0000006a;
			308: 	div_val = 32'h0000006a;
			309: 	div_val = 32'h0000006a;
			310: 	div_val = 32'h00000069;
			311: 	div_val = 32'h00000069;
			312: 	div_val = 32'h00000069;
			313: 	div_val = 32'h00000068;
			314: 	div_val = 32'h00000068;
			315: 	div_val = 32'h00000068;
			316: 	div_val = 32'h00000067;
			317: 	div_val = 32'h00000067;
			318: 	div_val = 32'h00000067;
			319: 	div_val = 32'h00000066;
			320: 	div_val = 32'h00000066;
			321: 	div_val = 32'h00000066;
			322: 	div_val = 32'h00000065;
			323: 	div_val = 32'h00000065;
			324: 	div_val = 32'h00000065;
			325: 	div_val = 32'h00000064;
			326: 	div_val = 32'h00000064;
			327: 	div_val = 32'h00000064;
			328: 	div_val = 32'h00000063;
			329: 	div_val = 32'h00000063;
			330: 	div_val = 32'h00000063;
			331: 	div_val = 32'h00000062;
			332: 	div_val = 32'h00000062;
			333: 	div_val = 32'h00000062;
			334: 	div_val = 32'h00000062;
			335: 	div_val = 32'h00000061;
			336: 	div_val = 32'h00000061;
			337: 	div_val = 32'h00000061;
			338: 	div_val = 32'h00000060;
			339: 	div_val = 32'h00000060;
			340: 	div_val = 32'h00000060;
			341: 	div_val = 32'h00000060;
			342: 	div_val = 32'h0000005f;
			343: 	div_val = 32'h0000005f;
			344: 	div_val = 32'h0000005f;
			345: 	div_val = 32'h0000005e;
			346: 	div_val = 32'h0000005e;
			347: 	div_val = 32'h0000005e;
			348: 	div_val = 32'h0000005e;
			349: 	div_val = 32'h0000005d;
			350: 	div_val = 32'h0000005d;
			351: 	div_val = 32'h0000005d;
			352: 	div_val = 32'h0000005d;
			353: 	div_val = 32'h0000005c;
			354: 	div_val = 32'h0000005c;
			355: 	div_val = 32'h0000005c;
			356: 	div_val = 32'h0000005c;
			357: 	div_val = 32'h0000005b;
			358: 	div_val = 32'h0000005b;
			359: 	div_val = 32'h0000005b;
			360: 	div_val = 32'h0000005b;
			361: 	div_val = 32'h0000005a;
			362: 	div_val = 32'h0000005a;
			363: 	div_val = 32'h0000005a;
			364: 	div_val = 32'h0000005a;
			365: 	div_val = 32'h00000059;
			366: 	div_val = 32'h00000059;
			367: 	div_val = 32'h00000059;
			368: 	div_val = 32'h00000059;
			369: 	div_val = 32'h00000058;
			370: 	div_val = 32'h00000058;
			371: 	div_val = 32'h00000058;
			372: 	div_val = 32'h00000058;
			373: 	div_val = 32'h00000057;
			374: 	div_val = 32'h00000057;
			375: 	div_val = 32'h00000057;
			376: 	div_val = 32'h00000057;
			377: 	div_val = 32'h00000056;
			378: 	div_val = 32'h00000056;
			379: 	div_val = 32'h00000056;
			380: 	div_val = 32'h00000056;
			381: 	div_val = 32'h00000056;
			382: 	div_val = 32'h00000055;
			383: 	div_val = 32'h00000055;
			384: 	div_val = 32'h00000055;
			385: 	div_val = 32'h00000055;
			386: 	div_val = 32'h00000054;
			387: 	div_val = 32'h00000054;
			388: 	div_val = 32'h00000054;
			389: 	div_val = 32'h00000054;
			390: 	div_val = 32'h00000054;
			391: 	div_val = 32'h00000053;
			392: 	div_val = 32'h00000053;
			393: 	div_val = 32'h00000053;
			394: 	div_val = 32'h00000053;
			395: 	div_val = 32'h00000052;
			396: 	div_val = 32'h00000052;
			397: 	div_val = 32'h00000052;
			398: 	div_val = 32'h00000052;
			399: 	div_val = 32'h00000052;
			400: 	div_val = 32'h00000051;
			401: 	div_val = 32'h00000051;
			402: 	div_val = 32'h00000051;
			403: 	div_val = 32'h00000051;
			404: 	div_val = 32'h00000051;
			405: 	div_val = 32'h00000050;
			406: 	div_val = 32'h00000050;
			407: 	div_val = 32'h00000050;
			408: 	div_val = 32'h00000050;
			409: 	div_val = 32'h00000050;
			410: 	div_val = 32'h0000004f;
			411: 	div_val = 32'h0000004f;
			412: 	div_val = 32'h0000004f;
			413: 	div_val = 32'h0000004f;
			414: 	div_val = 32'h0000004f;
			415: 	div_val = 32'h0000004e;
			416: 	div_val = 32'h0000004e;
			417: 	div_val = 32'h0000004e;
			418: 	div_val = 32'h0000004e;
			419: 	div_val = 32'h0000004e;
			420: 	div_val = 32'h0000004e;
			421: 	div_val = 32'h0000004d;
			422: 	div_val = 32'h0000004d;
			423: 	div_val = 32'h0000004d;
			424: 	div_val = 32'h0000004d;
			425: 	div_val = 32'h0000004d;
			426: 	div_val = 32'h0000004c;
			427: 	div_val = 32'h0000004c;
			428: 	div_val = 32'h0000004c;
			429: 	div_val = 32'h0000004c;
			430: 	div_val = 32'h0000004c;
			431: 	div_val = 32'h0000004c;
			432: 	div_val = 32'h0000004b;
			433: 	div_val = 32'h0000004b;
			434: 	div_val = 32'h0000004b;
			435: 	div_val = 32'h0000004b;
			436: 	div_val = 32'h0000004b;
			437: 	div_val = 32'h0000004a;
			438: 	div_val = 32'h0000004a;
			439: 	div_val = 32'h0000004a;
			440: 	div_val = 32'h0000004a;
			441: 	div_val = 32'h0000004a;
			442: 	div_val = 32'h0000004a;
			443: 	div_val = 32'h00000049;
			444: 	div_val = 32'h00000049;
			445: 	div_val = 32'h00000049;
			446: 	div_val = 32'h00000049;
			447: 	div_val = 32'h00000049;
			448: 	div_val = 32'h00000049;
			449: 	div_val = 32'h00000048;
			450: 	div_val = 32'h00000048;
			451: 	div_val = 32'h00000048;
			452: 	div_val = 32'h00000048;
			453: 	div_val = 32'h00000048;
			454: 	div_val = 32'h00000048;
			455: 	div_val = 32'h00000048;
			456: 	div_val = 32'h00000047;
			457: 	div_val = 32'h00000047;
			458: 	div_val = 32'h00000047;
			459: 	div_val = 32'h00000047;
			460: 	div_val = 32'h00000047;
			461: 	div_val = 32'h00000047;
			462: 	div_val = 32'h00000046;
			463: 	div_val = 32'h00000046;
			464: 	div_val = 32'h00000046;
			465: 	div_val = 32'h00000046;
			466: 	div_val = 32'h00000046;
			467: 	div_val = 32'h00000046;
			468: 	div_val = 32'h00000046;
			469: 	div_val = 32'h00000045;
			470: 	div_val = 32'h00000045;
			471: 	div_val = 32'h00000045;
			472: 	div_val = 32'h00000045;
			473: 	div_val = 32'h00000045;
			474: 	div_val = 32'h00000045;
			475: 	div_val = 32'h00000044;
			476: 	div_val = 32'h00000044;
			477: 	div_val = 32'h00000044;
			478: 	div_val = 32'h00000044;
			479: 	div_val = 32'h00000044;
			480: 	div_val = 32'h00000044;
			481: 	div_val = 32'h00000044;
			482: 	div_val = 32'h00000043;
			483: 	div_val = 32'h00000043;
			484: 	div_val = 32'h00000043;
			485: 	div_val = 32'h00000043;
			486: 	div_val = 32'h00000043;
			487: 	div_val = 32'h00000043;
			488: 	div_val = 32'h00000043;
			489: 	div_val = 32'h00000043;
			490: 	div_val = 32'h00000042;
			491: 	div_val = 32'h00000042;
			492: 	div_val = 32'h00000042;
			493: 	div_val = 32'h00000042;
			494: 	div_val = 32'h00000042;
			495: 	div_val = 32'h00000042;
			496: 	div_val = 32'h00000042;
			497: 	div_val = 32'h00000041;
			498: 	div_val = 32'h00000041;
			499: 	div_val = 32'h00000041;
			500: 	div_val = 32'h00000041;
			501: 	div_val = 32'h00000041;
			502: 	div_val = 32'h00000041;
			503: 	div_val = 32'h00000041;
			504: 	div_val = 32'h00000041;
			505: 	div_val = 32'h00000040;
			506: 	div_val = 32'h00000040;
			507: 	div_val = 32'h00000040;
			508: 	div_val = 32'h00000040;
			509: 	div_val = 32'h00000040;
			510: 	div_val = 32'h00000040;
			511: 	div_val = 32'h00000040;
			512: 	div_val = 32'h00000040;
			513: 	div_val = 32'h0000003f;
			514: 	div_val = 32'h0000003f;
			515: 	div_val = 32'h0000003f;
			516: 	div_val = 32'h0000003f;
			517: 	div_val = 32'h0000003f;
			518: 	div_val = 32'h0000003f;
			519: 	div_val = 32'h0000003f;
			520: 	div_val = 32'h0000003f;
			521: 	div_val = 32'h0000003e;
			522: 	div_val = 32'h0000003e;
			523: 	div_val = 32'h0000003e;
			524: 	div_val = 32'h0000003e;
			525: 	div_val = 32'h0000003e;
			526: 	div_val = 32'h0000003e;
			527: 	div_val = 32'h0000003e;
			528: 	div_val = 32'h0000003e;
			529: 	div_val = 32'h0000003d;
			530: 	div_val = 32'h0000003d;
			531: 	div_val = 32'h0000003d;
			532: 	div_val = 32'h0000003d;
			533: 	div_val = 32'h0000003d;
			534: 	div_val = 32'h0000003d;
			535: 	div_val = 32'h0000003d;
			536: 	div_val = 32'h0000003d;
			537: 	div_val = 32'h0000003d;
			538: 	div_val = 32'h0000003c;
			539: 	div_val = 32'h0000003c;
			540: 	div_val = 32'h0000003c;
			541: 	div_val = 32'h0000003c;
			542: 	div_val = 32'h0000003c;
			543: 	div_val = 32'h0000003c;
			544: 	div_val = 32'h0000003c;
			545: 	div_val = 32'h0000003c;
			546: 	div_val = 32'h0000003c;
			547: 	div_val = 32'h0000003b;
			548: 	div_val = 32'h0000003b;
			549: 	div_val = 32'h0000003b;
			550: 	div_val = 32'h0000003b;
			551: 	div_val = 32'h0000003b;
			552: 	div_val = 32'h0000003b;
			553: 	div_val = 32'h0000003b;
			554: 	div_val = 32'h0000003b;
			555: 	div_val = 32'h0000003b;
			556: 	div_val = 32'h0000003a;
			557: 	div_val = 32'h0000003a;
			558: 	div_val = 32'h0000003a;
			559: 	div_val = 32'h0000003a;
			560: 	div_val = 32'h0000003a;
			561: 	div_val = 32'h0000003a;
			562: 	div_val = 32'h0000003a;
			563: 	div_val = 32'h0000003a;
			564: 	div_val = 32'h0000003a;
			565: 	div_val = 32'h00000039;
			566: 	div_val = 32'h00000039;
			567: 	div_val = 32'h00000039;
			568: 	div_val = 32'h00000039;
			569: 	div_val = 32'h00000039;
			570: 	div_val = 32'h00000039;
			571: 	div_val = 32'h00000039;
			572: 	div_val = 32'h00000039;
			573: 	div_val = 32'h00000039;
			574: 	div_val = 32'h00000039;
			575: 	div_val = 32'h00000038;
			576: 	div_val = 32'h00000038;
			577: 	div_val = 32'h00000038;
			578: 	div_val = 32'h00000038;
			579: 	div_val = 32'h00000038;
			580: 	div_val = 32'h00000038;
			581: 	div_val = 32'h00000038;
			582: 	div_val = 32'h00000038;
			583: 	div_val = 32'h00000038;
			584: 	div_val = 32'h00000038;
			585: 	div_val = 32'h00000038;
			586: 	div_val = 32'h00000037;
			587: 	div_val = 32'h00000037;
			588: 	div_val = 32'h00000037;
			589: 	div_val = 32'h00000037;
			590: 	div_val = 32'h00000037;
			591: 	div_val = 32'h00000037;
			592: 	div_val = 32'h00000037;
			593: 	div_val = 32'h00000037;
			594: 	div_val = 32'h00000037;
			595: 	div_val = 32'h00000037;
			596: 	div_val = 32'h00000036;
			597: 	div_val = 32'h00000036;
			598: 	div_val = 32'h00000036;
			599: 	div_val = 32'h00000036;
			600: 	div_val = 32'h00000036;
			601: 	div_val = 32'h00000036;
			602: 	div_val = 32'h00000036;
			603: 	div_val = 32'h00000036;
			604: 	div_val = 32'h00000036;
			605: 	div_val = 32'h00000036;
			606: 	div_val = 32'h00000036;
			607: 	div_val = 32'h00000035;
			608: 	div_val = 32'h00000035;
			609: 	div_val = 32'h00000035;
			610: 	div_val = 32'h00000035;
			611: 	div_val = 32'h00000035;
			612: 	div_val = 32'h00000035;
			613: 	div_val = 32'h00000035;
			614: 	div_val = 32'h00000035;
			615: 	div_val = 32'h00000035;
			616: 	div_val = 32'h00000035;
			617: 	div_val = 32'h00000035;
			618: 	div_val = 32'h00000035;
			619: 	div_val = 32'h00000034;
			620: 	div_val = 32'h00000034;
			621: 	div_val = 32'h00000034;
			622: 	div_val = 32'h00000034;
			623: 	div_val = 32'h00000034;
			624: 	div_val = 32'h00000034;
			625: 	div_val = 32'h00000034;
			626: 	div_val = 32'h00000034;
			627: 	div_val = 32'h00000034;
			628: 	div_val = 32'h00000034;
			629: 	div_val = 32'h00000034;
			630: 	div_val = 32'h00000034;
			631: 	div_val = 32'h00000033;
			632: 	div_val = 32'h00000033;
			633: 	div_val = 32'h00000033;
			634: 	div_val = 32'h00000033;
			635: 	div_val = 32'h00000033;
			636: 	div_val = 32'h00000033;
			637: 	div_val = 32'h00000033;
			638: 	div_val = 32'h00000033;
			639: 	div_val = 32'h00000033;
			640: 	div_val = 32'h00000033;
			641: 	div_val = 32'h00000033;
			642: 	div_val = 32'h00000033;
			643: 	div_val = 32'h00000032;
			644: 	div_val = 32'h00000032;
			645: 	div_val = 32'h00000032;
			646: 	div_val = 32'h00000032;
			647: 	div_val = 32'h00000032;
			648: 	div_val = 32'h00000032;
			649: 	div_val = 32'h00000032;
			650: 	div_val = 32'h00000032;
			651: 	div_val = 32'h00000032;
			652: 	div_val = 32'h00000032;
			653: 	div_val = 32'h00000032;
			654: 	div_val = 32'h00000032;
			655: 	div_val = 32'h00000032;
			656: 	div_val = 32'h00000031;
			657: 	div_val = 32'h00000031;
			658: 	div_val = 32'h00000031;
			659: 	div_val = 32'h00000031;
			660: 	div_val = 32'h00000031;
			661: 	div_val = 32'h00000031;
			662: 	div_val = 32'h00000031;
			663: 	div_val = 32'h00000031;
			664: 	div_val = 32'h00000031;
			665: 	div_val = 32'h00000031;
			666: 	div_val = 32'h00000031;
			667: 	div_val = 32'h00000031;
			668: 	div_val = 32'h00000031;
			669: 	div_val = 32'h00000030;
			670: 	div_val = 32'h00000030;
			671: 	div_val = 32'h00000030;
			672: 	div_val = 32'h00000030;
			673: 	div_val = 32'h00000030;
			674: 	div_val = 32'h00000030;
			675: 	div_val = 32'h00000030;
			676: 	div_val = 32'h00000030;
			677: 	div_val = 32'h00000030;
			678: 	div_val = 32'h00000030;
			679: 	div_val = 32'h00000030;
			680: 	div_val = 32'h00000030;
			681: 	div_val = 32'h00000030;
			682: 	div_val = 32'h00000030;
			683: 	div_val = 32'h0000002f;
			684: 	div_val = 32'h0000002f;
			685: 	div_val = 32'h0000002f;
			686: 	div_val = 32'h0000002f;
			687: 	div_val = 32'h0000002f;
			688: 	div_val = 32'h0000002f;
			689: 	div_val = 32'h0000002f;
			690: 	div_val = 32'h0000002f;
			691: 	div_val = 32'h0000002f;
			692: 	div_val = 32'h0000002f;
			693: 	div_val = 32'h0000002f;
			694: 	div_val = 32'h0000002f;
			695: 	div_val = 32'h0000002f;
			696: 	div_val = 32'h0000002f;
			697: 	div_val = 32'h0000002f;
			698: 	div_val = 32'h0000002e;
			699: 	div_val = 32'h0000002e;
			700: 	div_val = 32'h0000002e;
			701: 	div_val = 32'h0000002e;
			702: 	div_val = 32'h0000002e;
			703: 	div_val = 32'h0000002e;
			704: 	div_val = 32'h0000002e;
			705: 	div_val = 32'h0000002e;
			706: 	div_val = 32'h0000002e;
			707: 	div_val = 32'h0000002e;
			708: 	div_val = 32'h0000002e;
			709: 	div_val = 32'h0000002e;
			710: 	div_val = 32'h0000002e;
			711: 	div_val = 32'h0000002e;
			712: 	div_val = 32'h0000002e;
			713: 	div_val = 32'h0000002d;
			714: 	div_val = 32'h0000002d;
			715: 	div_val = 32'h0000002d;
			716: 	div_val = 32'h0000002d;
			717: 	div_val = 32'h0000002d;
			718: 	div_val = 32'h0000002d;
			719: 	div_val = 32'h0000002d;
			720: 	div_val = 32'h0000002d;
			721: 	div_val = 32'h0000002d;
			722: 	div_val = 32'h0000002d;
			723: 	div_val = 32'h0000002d;
			724: 	div_val = 32'h0000002d;
			725: 	div_val = 32'h0000002d;
			726: 	div_val = 32'h0000002d;
			727: 	div_val = 32'h0000002d;
			728: 	div_val = 32'h0000002d;
			729: 	div_val = 32'h0000002c;
			730: 	div_val = 32'h0000002c;
			731: 	div_val = 32'h0000002c;
			732: 	div_val = 32'h0000002c;
			733: 	div_val = 32'h0000002c;
			734: 	div_val = 32'h0000002c;
			735: 	div_val = 32'h0000002c;
			736: 	div_val = 32'h0000002c;
			737: 	div_val = 32'h0000002c;
			738: 	div_val = 32'h0000002c;
			739: 	div_val = 32'h0000002c;
			740: 	div_val = 32'h0000002c;
			741: 	div_val = 32'h0000002c;
			742: 	div_val = 32'h0000002c;
			743: 	div_val = 32'h0000002c;
			744: 	div_val = 32'h0000002c;
			745: 	div_val = 32'h0000002b;
			746: 	div_val = 32'h0000002b;
			747: 	div_val = 32'h0000002b;
			748: 	div_val = 32'h0000002b;
			749: 	div_val = 32'h0000002b;
			750: 	div_val = 32'h0000002b;
			751: 	div_val = 32'h0000002b;
			752: 	div_val = 32'h0000002b;
			753: 	div_val = 32'h0000002b;
			754: 	div_val = 32'h0000002b;
			755: 	div_val = 32'h0000002b;
			756: 	div_val = 32'h0000002b;
			757: 	div_val = 32'h0000002b;
			758: 	div_val = 32'h0000002b;
			759: 	div_val = 32'h0000002b;
			760: 	div_val = 32'h0000002b;
			761: 	div_val = 32'h0000002b;
			762: 	div_val = 32'h0000002b;
			763: 	div_val = 32'h0000002a;
			764: 	div_val = 32'h0000002a;
			765: 	div_val = 32'h0000002a;
			766: 	div_val = 32'h0000002a;
			767: 	div_val = 32'h0000002a;
			768: 	div_val = 32'h0000002a;
			769: 	div_val = 32'h0000002a;
			770: 	div_val = 32'h0000002a;
			771: 	div_val = 32'h0000002a;
			772: 	div_val = 32'h0000002a;
			773: 	div_val = 32'h0000002a;
			774: 	div_val = 32'h0000002a;
			775: 	div_val = 32'h0000002a;
			776: 	div_val = 32'h0000002a;
			777: 	div_val = 32'h0000002a;
			778: 	div_val = 32'h0000002a;
			779: 	div_val = 32'h0000002a;
			780: 	div_val = 32'h0000002a;
			781: 	div_val = 32'h00000029;
			782: 	div_val = 32'h00000029;
			783: 	div_val = 32'h00000029;
			784: 	div_val = 32'h00000029;
			785: 	div_val = 32'h00000029;
			786: 	div_val = 32'h00000029;
			787: 	div_val = 32'h00000029;
			788: 	div_val = 32'h00000029;
			789: 	div_val = 32'h00000029;
			790: 	div_val = 32'h00000029;
			791: 	div_val = 32'h00000029;
			792: 	div_val = 32'h00000029;
			793: 	div_val = 32'h00000029;
			794: 	div_val = 32'h00000029;
			795: 	div_val = 32'h00000029;
			796: 	div_val = 32'h00000029;
			797: 	div_val = 32'h00000029;
			798: 	div_val = 32'h00000029;
			799: 	div_val = 32'h00000029;
			800: 	div_val = 32'h00000028;
			801: 	div_val = 32'h00000028;
			802: 	div_val = 32'h00000028;
			803: 	div_val = 32'h00000028;
			804: 	div_val = 32'h00000028;
			805: 	div_val = 32'h00000028;
			806: 	div_val = 32'h00000028;
			807: 	div_val = 32'h00000028;
			808: 	div_val = 32'h00000028;
			809: 	div_val = 32'h00000028;
			810: 	div_val = 32'h00000028;
			811: 	div_val = 32'h00000028;
			812: 	div_val = 32'h00000028;
			813: 	div_val = 32'h00000028;
			814: 	div_val = 32'h00000028;
			815: 	div_val = 32'h00000028;
			816: 	div_val = 32'h00000028;
			817: 	div_val = 32'h00000028;
			818: 	div_val = 32'h00000028;
			819: 	div_val = 32'h00000028;
			820: 	div_val = 32'h00000027;
			821: 	div_val = 32'h00000027;
			822: 	div_val = 32'h00000027;
			823: 	div_val = 32'h00000027;
			824: 	div_val = 32'h00000027;
			825: 	div_val = 32'h00000027;
			826: 	div_val = 32'h00000027;
			827: 	div_val = 32'h00000027;
			828: 	div_val = 32'h00000027;
			829: 	div_val = 32'h00000027;
			830: 	div_val = 32'h00000027;
			831: 	div_val = 32'h00000027;
			832: 	div_val = 32'h00000027;
			833: 	div_val = 32'h00000027;
			834: 	div_val = 32'h00000027;
			835: 	div_val = 32'h00000027;
			836: 	div_val = 32'h00000027;
			837: 	div_val = 32'h00000027;
			838: 	div_val = 32'h00000027;
			839: 	div_val = 32'h00000027;
			840: 	div_val = 32'h00000027;
			841: 	div_val = 32'h00000026;
			842: 	div_val = 32'h00000026;
			843: 	div_val = 32'h00000026;
			844: 	div_val = 32'h00000026;
			845: 	div_val = 32'h00000026;
			846: 	div_val = 32'h00000026;
			847: 	div_val = 32'h00000026;
			848: 	div_val = 32'h00000026;
			849: 	div_val = 32'h00000026;
			850: 	div_val = 32'h00000026;
			851: 	div_val = 32'h00000026;
			852: 	div_val = 32'h00000026;
			853: 	div_val = 32'h00000026;
			854: 	div_val = 32'h00000026;
			855: 	div_val = 32'h00000026;
			856: 	div_val = 32'h00000026;
			857: 	div_val = 32'h00000026;
			858: 	div_val = 32'h00000026;
			859: 	div_val = 32'h00000026;
			860: 	div_val = 32'h00000026;
			861: 	div_val = 32'h00000026;
			862: 	div_val = 32'h00000026;
			863: 	div_val = 32'h00000025;
			864: 	div_val = 32'h00000025;
			865: 	div_val = 32'h00000025;
			866: 	div_val = 32'h00000025;
			867: 	div_val = 32'h00000025;
			868: 	div_val = 32'h00000025;
			869: 	div_val = 32'h00000025;
			870: 	div_val = 32'h00000025;
			871: 	div_val = 32'h00000025;
			872: 	div_val = 32'h00000025;
			873: 	div_val = 32'h00000025;
			874: 	div_val = 32'h00000025;
			875: 	div_val = 32'h00000025;
			876: 	div_val = 32'h00000025;
			877: 	div_val = 32'h00000025;
			878: 	div_val = 32'h00000025;
			879: 	div_val = 32'h00000025;
			880: 	div_val = 32'h00000025;
			881: 	div_val = 32'h00000025;
			882: 	div_val = 32'h00000025;
			883: 	div_val = 32'h00000025;
			884: 	div_val = 32'h00000025;
			885: 	div_val = 32'h00000025;
			886: 	div_val = 32'h00000024;
			887: 	div_val = 32'h00000024;
			888: 	div_val = 32'h00000024;
			889: 	div_val = 32'h00000024;
			890: 	div_val = 32'h00000024;
			891: 	div_val = 32'h00000024;
			892: 	div_val = 32'h00000024;
			893: 	div_val = 32'h00000024;
			894: 	div_val = 32'h00000024;
			895: 	div_val = 32'h00000024;
			896: 	div_val = 32'h00000024;
			897: 	div_val = 32'h00000024;
			898: 	div_val = 32'h00000024;
			899: 	div_val = 32'h00000024;
			900: 	div_val = 32'h00000024;
			901: 	div_val = 32'h00000024;
			902: 	div_val = 32'h00000024;
			903: 	div_val = 32'h00000024;
			904: 	div_val = 32'h00000024;
			905: 	div_val = 32'h00000024;
			906: 	div_val = 32'h00000024;
			907: 	div_val = 32'h00000024;
			908: 	div_val = 32'h00000024;
			909: 	div_val = 32'h00000024;
			910: 	div_val = 32'h00000024;
			911: 	div_val = 32'h00000023;
			912: 	div_val = 32'h00000023;
			913: 	div_val = 32'h00000023;
			914: 	div_val = 32'h00000023;
			915: 	div_val = 32'h00000023;
			916: 	div_val = 32'h00000023;
			917: 	div_val = 32'h00000023;
			918: 	div_val = 32'h00000023;
			919: 	div_val = 32'h00000023;
			920: 	div_val = 32'h00000023;
			921: 	div_val = 32'h00000023;
			922: 	div_val = 32'h00000023;
			923: 	div_val = 32'h00000023;
			924: 	div_val = 32'h00000023;
			925: 	div_val = 32'h00000023;
			926: 	div_val = 32'h00000023;
			927: 	div_val = 32'h00000023;
			928: 	div_val = 32'h00000023;
			929: 	div_val = 32'h00000023;
			930: 	div_val = 32'h00000023;
			931: 	div_val = 32'h00000023;
			932: 	div_val = 32'h00000023;
			933: 	div_val = 32'h00000023;
			934: 	div_val = 32'h00000023;
			935: 	div_val = 32'h00000023;
			936: 	div_val = 32'h00000023;
			937: 	div_val = 32'h00000022;
			938: 	div_val = 32'h00000022;
			939: 	div_val = 32'h00000022;
			940: 	div_val = 32'h00000022;
			941: 	div_val = 32'h00000022;
			942: 	div_val = 32'h00000022;
			943: 	div_val = 32'h00000022;
			944: 	div_val = 32'h00000022;
			945: 	div_val = 32'h00000022;
			946: 	div_val = 32'h00000022;
			947: 	div_val = 32'h00000022;
			948: 	div_val = 32'h00000022;
			949: 	div_val = 32'h00000022;
			950: 	div_val = 32'h00000022;
			951: 	div_val = 32'h00000022;
			952: 	div_val = 32'h00000022;
			953: 	div_val = 32'h00000022;
			954: 	div_val = 32'h00000022;
			955: 	div_val = 32'h00000022;
			956: 	div_val = 32'h00000022;
			957: 	div_val = 32'h00000022;
			958: 	div_val = 32'h00000022;
			959: 	div_val = 32'h00000022;
			960: 	div_val = 32'h00000022;
			961: 	div_val = 32'h00000022;
			962: 	div_val = 32'h00000022;
			963: 	div_val = 32'h00000022;
			964: 	div_val = 32'h00000021;
			965: 	div_val = 32'h00000021;
			966: 	div_val = 32'h00000021;
			967: 	div_val = 32'h00000021;
			968: 	div_val = 32'h00000021;
			969: 	div_val = 32'h00000021;
			970: 	div_val = 32'h00000021;
			971: 	div_val = 32'h00000021;
			972: 	div_val = 32'h00000021;
			973: 	div_val = 32'h00000021;
			974: 	div_val = 32'h00000021;
			975: 	div_val = 32'h00000021;
			976: 	div_val = 32'h00000021;
			977: 	div_val = 32'h00000021;
			978: 	div_val = 32'h00000021;
			979: 	div_val = 32'h00000021;
			980: 	div_val = 32'h00000021;
			981: 	div_val = 32'h00000021;
			982: 	div_val = 32'h00000021;
			983: 	div_val = 32'h00000021;
			984: 	div_val = 32'h00000021;
			985: 	div_val = 32'h00000021;
			986: 	div_val = 32'h00000021;
			987: 	div_val = 32'h00000021;
			988: 	div_val = 32'h00000021;
			989: 	div_val = 32'h00000021;
			990: 	div_val = 32'h00000021;
			991: 	div_val = 32'h00000021;
			992: 	div_val = 32'h00000021;
			993: 	div_val = 32'h00000020;
			994: 	div_val = 32'h00000020;
			995: 	div_val = 32'h00000020;
			996: 	div_val = 32'h00000020;
			997: 	div_val = 32'h00000020;
			998: 	div_val = 32'h00000020;
			999: 	div_val = 32'h00000020;
			1000: 	div_val = 32'h00000020;
			1001: 	div_val = 32'h00000020;
			1002: 	div_val = 32'h00000020;
			1003: 	div_val = 32'h00000020;
			1004: 	div_val = 32'h00000020;
			1005: 	div_val = 32'h00000020;
			1006: 	div_val = 32'h00000020;
			1007: 	div_val = 32'h00000020;
			1008: 	div_val = 32'h00000020;
			1009: 	div_val = 32'h00000020;
			1010: 	div_val = 32'h00000020;
			1011: 	div_val = 32'h00000020;
			1012: 	div_val = 32'h00000020;
			1013: 	div_val = 32'h00000020;
			1014: 	div_val = 32'h00000020;
			1015: 	div_val = 32'h00000020;
			1016: 	div_val = 32'h00000020;
			1017: 	div_val = 32'h00000020;
			1018: 	div_val = 32'h00000020;
			1019: 	div_val = 32'h00000020;
			1020: 	div_val = 32'h00000020;
			1021: 	div_val = 32'h00000020;
			1022: 	div_val = 32'h00000020;
			1023: 	div_val = 32'h00000020;
			default: div_val = 32'b0;
		endcase
	end

endmodule